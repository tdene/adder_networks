
module adder(cout, sum, a, b, cin);
	input [31:0] a, b;
	input cin;
	output [31:0] sum;
	output cout;
	wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, g_lsb, p_lsb, g0, p0, g1, p1, g2, p2, g3, p3, g4, p4, g5, p5, g6, p6, g7, p7, g8, p8, g9, p9, g10, p10, g11, p11, g12, p12, g13, p13, g14, p14, g15, p15, g16, p16, g17, p17, g18, p18, g19, p19, g20, p20, g21, p21, g22, p22, g23, p23, g24, p24, g25, p25, g26, p26, g27, p27, g28, p28, g29, p29, g30, p30, g31, p31;
	pre_node pre_node_32_0 ( .a_in( a[31] ), .b_in( b[31] ), .pout ( p31 ), .gout ( g31 ) );
	grey grey_node_cout ( .gin ( {g31,n544} ), .pin ( p31 ), .gout ( cout ) );
	fake_pre fake_pre_0_0 ( .cin( {cin} ), .pout( {p_lsb} ), .gout( {g_lsb} ) );
	pre_node pre_node_1_0 ( .a_in( {a[0]} ), .b_in( {b[0]} ), .pout( {p0} ), .gout( {g0} ) );
	pre_node pre_node_2_0 ( .a_in( {a[1]} ), .b_in( {b[1]} ), .pout( {p1} ), .gout( {g1} ) );
	pre_node pre_node_3_0 ( .a_in( {a[2]} ), .b_in( {b[2]} ), .pout( {p2} ), .gout( {g2} ) );
	pre_node pre_node_4_0 ( .a_in( {a[3]} ), .b_in( {b[3]} ), .pout( {p3} ), .gout( {g3} ) );
	pre_node pre_node_5_0 ( .a_in( {a[4]} ), .b_in( {b[4]} ), .pout( {p4} ), .gout( {g4} ) );
	pre_node pre_node_6_0 ( .a_in( {a[5]} ), .b_in( {b[5]} ), .pout( {p5} ), .gout( {g5} ) );
	pre_node pre_node_7_0 ( .a_in( {a[6]} ), .b_in( {b[6]} ), .pout( {p6} ), .gout( {g6} ) );
	pre_node pre_node_8_0 ( .a_in( {a[7]} ), .b_in( {b[7]} ), .pout( {p7} ), .gout( {g7} ) );
	pre_node pre_node_9_0 ( .a_in( {a[8]} ), .b_in( {b[8]} ), .pout( {p8} ), .gout( {g8} ) );
	pre_node pre_node_10_0 ( .a_in( {a[9]} ), .b_in( {b[9]} ), .pout( {p9} ), .gout( {g9} ) );
	pre_node pre_node_11_0 ( .a_in( {a[10]} ), .b_in( {b[10]} ), .pout( {p10} ), .gout( {g10} ) );
	pre_node pre_node_12_0 ( .a_in( {a[11]} ), .b_in( {b[11]} ), .pout( {p11} ), .gout( {g11} ) );
	pre_node pre_node_13_0 ( .a_in( {a[12]} ), .b_in( {b[12]} ), .pout( {p12} ), .gout( {g12} ) );
	pre_node pre_node_14_0 ( .a_in( {a[13]} ), .b_in( {b[13]} ), .pout( {p13} ), .gout( {g13} ) );
	pre_node pre_node_15_0 ( .a_in( {a[14]} ), .b_in( {b[14]} ), .pout( {p14} ), .gout( {g14} ) );
	pre_node pre_node_16_0 ( .a_in( {a[15]} ), .b_in( {b[15]} ), .pout( {p15} ), .gout( {g15} ) );
	pre_node pre_node_17_0 ( .a_in( {a[16]} ), .b_in( {b[16]} ), .pout( {p16} ), .gout( {g16} ) );
	pre_node pre_node_18_0 ( .a_in( {a[17]} ), .b_in( {b[17]} ), .pout( {p17} ), .gout( {g17} ) );
	pre_node pre_node_19_0 ( .a_in( {a[18]} ), .b_in( {b[18]} ), .pout( {p18} ), .gout( {g18} ) );
	pre_node pre_node_20_0 ( .a_in( {a[19]} ), .b_in( {b[19]} ), .pout( {p19} ), .gout( {g19} ) );
	pre_node pre_node_21_0 ( .a_in( {a[20]} ), .b_in( {b[20]} ), .pout( {p20} ), .gout( {g20} ) );
	pre_node pre_node_22_0 ( .a_in( {a[21]} ), .b_in( {b[21]} ), .pout( {p21} ), .gout( {g21} ) );
	pre_node pre_node_23_0 ( .a_in( {a[22]} ), .b_in( {b[22]} ), .pout( {p22} ), .gout( {g22} ) );
	pre_node pre_node_24_0 ( .a_in( {a[23]} ), .b_in( {b[23]} ), .pout( {p23} ), .gout( {g23} ) );
	pre_node pre_node_25_0 ( .a_in( {a[24]} ), .b_in( {b[24]} ), .pout( {p24} ), .gout( {g24} ) );
	pre_node pre_node_26_0 ( .a_in( {a[25]} ), .b_in( {b[25]} ), .pout( {p25} ), .gout( {g25} ) );
	pre_node pre_node_27_0 ( .a_in( {a[26]} ), .b_in( {b[26]} ), .pout( {p26} ), .gout( {g26} ) );
	pre_node pre_node_28_0 ( .a_in( {a[27]} ), .b_in( {b[27]} ), .pout( {p27} ), .gout( {g27} ) );
	pre_node pre_node_29_0 ( .a_in( {a[28]} ), .b_in( {b[28]} ), .pout( {p28} ), .gout( {g28} ) );
	pre_node pre_node_30_0 ( .a_in( {a[29]} ), .b_in( {b[29]} ), .pout( {p29} ), .gout( {g29} ) );
	pre_node pre_node_31_0 ( .a_in( {a[30]} ), .b_in( {b[30]} ), .pout( {p30} ), .gout( {g30} ) );
    assign n97=p_lsb;
    assign n98=g_lsb;

	black black_1_1 ( .gin( {g0,g_lsb} ), .pin( {p0,p_lsb} ), .gout( {n100} ), .pout( {n99} ) );
    assign n101=p1;
    assign n102=g1;

	black black_3_1 ( .gin( {g2,g1} ), .pin( {p2,p1} ), .gout( {n106} ), .pout( {n105} ) );
    assign n109=p3;
    assign n110=g3;

	black black_5_1 ( .gin( {g4,g3} ), .pin( {p4,p3} ), .gout( {n112} ), .pout( {n111} ) );
    assign n113=p5;
    assign n114=g5;

	black black_7_1 ( .gin( {g6,g5} ), .pin( {p6,p5} ), .gout( {n118} ), .pout( {n117} ) );
    assign n121=p7;
    assign n122=g7;

	black black_9_1 ( .gin( {g8,g7} ), .pin( {p8,p7} ), .gout( {n124} ), .pout( {n123} ) );
    assign n125=p9;
    assign n126=g9;

	black black_11_1 ( .gin( {g10,g9} ), .pin( {p10,p9} ), .gout( {n130} ), .pout( {n129} ) );
    assign n133=p11;
    assign n134=g11;

	black black_13_1 ( .gin( {g12,g11} ), .pin( {p12,p11} ), .gout( {n136} ), .pout( {n135} ) );
    assign n137=p13;
    assign n138=g13;

	black black_15_1 ( .gin( {g14,g13} ), .pin( {p14,p13} ), .gout( {n142} ), .pout( {n141} ) );
    assign n145=p15;
    assign n146=g15;

	black black_17_1 ( .gin( {g16,g15} ), .pin( {p16,p15} ), .gout( {n148} ), .pout( {n147} ) );
    assign n149=p17;
    assign n150=g17;

	black black_19_1 ( .gin( {g18,g17} ), .pin( {p18,p17} ), .gout( {n154} ), .pout( {n153} ) );
    assign n157=p19;
    assign n158=g19;

	black black_21_1 ( .gin( {g20,g19} ), .pin( {p20,p19} ), .gout( {n160} ), .pout( {n159} ) );
    assign n161=p21;
    assign n162=g21;

	black black_23_1 ( .gin( {g22,g21} ), .pin( {p22,p21} ), .gout( {n166} ), .pout( {n165} ) );
    assign n169=p23;
    assign n170=g23;

	black black_25_1 ( .gin( {g24,g23} ), .pin( {p24,p23} ), .gout( {n172} ), .pout( {n171} ) );
    assign n173=p25;
    assign n174=g25;

	black black_27_1 ( .gin( {g26,g25} ), .pin( {p26,p25} ), .gout( {n178} ), .pout( {n177} ) );
    assign n181=p27;
    assign n182=g27;

	black black_29_1 ( .gin( {g28,g27} ), .pin( {p28,p27} ), .gout( {n184} ), .pout( {n183} ) );
    assign n185=p29;
    assign n186=g29;

	black black_31_1 ( .gin( {g30,g29} ), .pin( {p30,p29} ), .gout( {n190} ), .pout( {n189} ) );
    assign n193=n97;
    assign n194=n98;

    assign n195=n99;
    assign n196=n100;

	black black_2_2 ( .gin( {n102,n100} ), .pin( {n101,n99} ), .gout( {n198} ), .pout( {n197} ) );
	black black_3_2 ( .gin( {n106,n100} ), .pin( {n105,n99} ), .gout( {n200} ), .pout( {n199} ) );
    assign n201=n109;
    assign n202=n110;

    assign n205=n111;
    assign n206=n112;

	black black_6_2 ( .gin( {n114,n112} ), .pin( {n113,n111} ), .gout( {n210} ), .pout( {n209} ) );
	black black_7_2 ( .gin( {n118,n112} ), .pin( {n117,n111} ), .gout( {n214} ), .pout( {n213} ) );
    assign n217=n121;
    assign n218=n122;

    assign n219=n123;
    assign n220=n124;

	black black_10_2 ( .gin( {n126,n124} ), .pin( {n125,n123} ), .gout( {n222} ), .pout( {n221} ) );
	black black_11_2 ( .gin( {n130,n124} ), .pin( {n129,n123} ), .gout( {n224} ), .pout( {n223} ) );
    assign n225=n133;
    assign n226=n134;

    assign n229=n135;
    assign n230=n136;

	black black_14_2 ( .gin( {n138,n136} ), .pin( {n137,n135} ), .gout( {n234} ), .pout( {n233} ) );
	black black_15_2 ( .gin( {n142,n136} ), .pin( {n141,n135} ), .gout( {n238} ), .pout( {n237} ) );
    assign n241=n145;
    assign n242=n146;

    assign n243=n147;
    assign n244=n148;

	black black_18_2 ( .gin( {n150,n148} ), .pin( {n149,n147} ), .gout( {n246} ), .pout( {n245} ) );
	black black_19_2 ( .gin( {n154,n148} ), .pin( {n153,n147} ), .gout( {n248} ), .pout( {n247} ) );
    assign n249=n157;
    assign n250=n158;

    assign n253=n159;
    assign n254=n160;

	black black_22_2 ( .gin( {n162,n160} ), .pin( {n161,n159} ), .gout( {n258} ), .pout( {n257} ) );
	black black_23_2 ( .gin( {n166,n160} ), .pin( {n165,n159} ), .gout( {n262} ), .pout( {n261} ) );
    assign n265=n169;
    assign n266=n170;

    assign n267=n171;
    assign n268=n172;

	black black_26_2 ( .gin( {n174,n172} ), .pin( {n173,n171} ), .gout( {n270} ), .pout( {n269} ) );
	black black_27_2 ( .gin( {n178,n172} ), .pin( {n177,n171} ), .gout( {n272} ), .pout( {n271} ) );
    assign n273=n181;
    assign n274=n182;

    assign n277=n183;
    assign n278=n184;

	black black_30_2 ( .gin( {n186,n184} ), .pin( {n185,n183} ), .gout( {n282} ), .pout( {n281} ) );
	black black_31_2 ( .gin( {n190,n184} ), .pin( {n189,n183} ), .gout( {n286} ), .pout( {n285} ) );
    assign n289=n193;
    assign n290=n194;

    assign n291=n195;
    assign n292=n196;

    assign n293=n197;
    assign n294=n198;

    assign n295=n199;
    assign n296=n200;

	black black_4_3 ( .gin( {n202,n200} ), .pin( {n201,n199} ), .gout( {n298} ), .pout( {n297} ) );
	black black_5_3 ( .gin( {n206,n200} ), .pin( {n205,n199} ), .gout( {n300} ), .pout( {n299} ) );
	black black_6_3 ( .gin( {n210,n200} ), .pin( {n209,n199} ), .gout( {n302} ), .pout( {n301} ) );
	black black_7_3 ( .gin( {n214,n200} ), .pin( {n213,n199} ), .gout( {n304} ), .pout( {n303} ) );
    assign n305=n217;
    assign n306=n218;

    assign n309=n219;
    assign n310=n220;

    assign n313=n221;
    assign n314=n222;

    assign n317=n223;
    assign n318=n224;

	black black_12_3 ( .gin( {n226,n224} ), .pin( {n225,n223} ), .gout( {n322} ), .pout( {n321} ) );
	black black_13_3 ( .gin( {n230,n224} ), .pin( {n229,n223} ), .gout( {n326} ), .pout( {n325} ) );
	black black_14_3 ( .gin( {n234,n224} ), .pin( {n233,n223} ), .gout( {n330} ), .pout( {n329} ) );
	black black_15_3 ( .gin( {n238,n224} ), .pin( {n237,n223} ), .gout( {n334} ), .pout( {n333} ) );
    assign n337=n241;
    assign n338=n242;

    assign n339=n243;
    assign n340=n244;

    assign n341=n245;
    assign n342=n246;

    assign n343=n247;
    assign n344=n248;

	black black_20_3 ( .gin( {n250,n248} ), .pin( {n249,n247} ), .gout( {n346} ), .pout( {n345} ) );
	black black_21_3 ( .gin( {n254,n248} ), .pin( {n253,n247} ), .gout( {n348} ), .pout( {n347} ) );
	black black_22_3 ( .gin( {n258,n248} ), .pin( {n257,n247} ), .gout( {n350} ), .pout( {n349} ) );
	black black_23_3 ( .gin( {n262,n248} ), .pin( {n261,n247} ), .gout( {n352} ), .pout( {n351} ) );
    assign n353=n265;
    assign n354=n266;

    assign n357=n267;
    assign n358=n268;

    assign n361=n269;
    assign n362=n270;

    assign n365=n271;
    assign n366=n272;

	black black_28_3 ( .gin( {n274,n272} ), .pin( {n273,n271} ), .gout( {n370} ), .pout( {n369} ) );
	black black_29_3 ( .gin( {n278,n272} ), .pin( {n277,n271} ), .gout( {n374} ), .pout( {n373} ) );
	black black_30_3 ( .gin( {n282,n272} ), .pin( {n281,n271} ), .gout( {n378} ), .pout( {n377} ) );
	black black_31_3 ( .gin( {n286,n272} ), .pin( {n285,n271} ), .gout( {n382} ), .pout( {n381} ) );
    assign n385=n289;
    assign n386=n290;

    assign n387=n291;
    assign n388=n292;

    assign n389=n293;
    assign n390=n294;

    assign n391=n295;
    assign n392=n296;

    assign n393=n297;
    assign n394=n298;

    assign n395=n299;
    assign n396=n300;

    assign n397=n301;
    assign n398=n302;

    assign n399=n303;
    assign n400=n304;

	black black_8_4 ( .gin( {n306,n304} ), .pin( {n305,n303} ), .gout( {n402} ), .pout( {n401} ) );
	black black_9_4 ( .gin( {n310,n304} ), .pin( {n309,n303} ), .gout( {n404} ), .pout( {n403} ) );
	black black_10_4 ( .gin( {n314,n304} ), .pin( {n313,n303} ), .gout( {n406} ), .pout( {n405} ) );
	black black_11_4 ( .gin( {n318,n304} ), .pin( {n317,n303} ), .gout( {n408} ), .pout( {n407} ) );
	black black_12_4 ( .gin( {n322,n304} ), .pin( {n321,n303} ), .gout( {n410} ), .pout( {n409} ) );
	black black_13_4 ( .gin( {n326,n304} ), .pin( {n325,n303} ), .gout( {n412} ), .pout( {n411} ) );
	black black_14_4 ( .gin( {n330,n304} ), .pin( {n329,n303} ), .gout( {n414} ), .pout( {n413} ) );
	black black_15_4 ( .gin( {n334,n304} ), .pin( {n333,n303} ), .gout( {n416} ), .pout( {n415} ) );
    assign n417=n337;
    assign n418=n338;

    assign n421=n339;
    assign n422=n340;

    assign n425=n341;
    assign n426=n342;

    assign n429=n343;
    assign n430=n344;

    assign n433=n345;
    assign n434=n346;

    assign n437=n347;
    assign n438=n348;

    assign n441=n349;
    assign n442=n350;

    assign n445=n351;
    assign n446=n352;

	black black_24_4 ( .gin( {n354,n352} ), .pin( {n353,n351} ), .gout( {n450} ), .pout( {n449} ) );
	black black_25_4 ( .gin( {n358,n352} ), .pin( {n357,n351} ), .gout( {n454} ), .pout( {n453} ) );
	black black_26_4 ( .gin( {n362,n352} ), .pin( {n361,n351} ), .gout( {n458} ), .pout( {n457} ) );
	black black_27_4 ( .gin( {n366,n352} ), .pin( {n365,n351} ), .gout( {n462} ), .pout( {n461} ) );
	black black_28_4 ( .gin( {n370,n352} ), .pin( {n369,n351} ), .gout( {n466} ), .pout( {n465} ) );
	black black_29_4 ( .gin( {n374,n352} ), .pin( {n373,n351} ), .gout( {n470} ), .pout( {n469} ) );
	black black_30_4 ( .gin( {n378,n352} ), .pin( {n377,n351} ), .gout( {n474} ), .pout( {n473} ) );
	black black_31_4 ( .gin( {n382,n352} ), .pin( {n381,n351} ), .gout( {n478} ), .pout( {n477} ) );
    assign n481=n385;
    assign n482=n386;

    assign n483=n387;
    assign n484=n388;

    assign n485=n389;
    assign n486=n390;

    assign n487=n391;
    assign n488=n392;

    assign n489=n393;
    assign n490=n394;

    assign n491=n395;
    assign n492=n396;

    assign n493=n397;
    assign n494=n398;

    assign n495=n399;
    assign n496=n400;

    assign n497=n401;
    assign n498=n402;

    assign n499=n403;
    assign n500=n404;

    assign n501=n405;
    assign n502=n406;

    assign n503=n407;
    assign n504=n408;

    assign n505=n409;
    assign n506=n410;

    assign n507=n411;
    assign n508=n412;

    assign n509=n413;
    assign n510=n414;

    assign n511=n415;
    assign n512=n416;

	black black_16_5 ( .gin( {n418,n416} ), .pin( {n417,n415} ), .gout( {n514} ), .pout( {n513} ) );
	black black_17_5 ( .gin( {n422,n416} ), .pin( {n421,n415} ), .gout( {n516} ), .pout( {n515} ) );
	black black_18_5 ( .gin( {n426,n416} ), .pin( {n425,n415} ), .gout( {n518} ), .pout( {n517} ) );
	black black_19_5 ( .gin( {n430,n416} ), .pin( {n429,n415} ), .gout( {n520} ), .pout( {n519} ) );
	black black_20_5 ( .gin( {n434,n416} ), .pin( {n433,n415} ), .gout( {n522} ), .pout( {n521} ) );
	black black_21_5 ( .gin( {n438,n416} ), .pin( {n437,n415} ), .gout( {n524} ), .pout( {n523} ) );
	black black_22_5 ( .gin( {n442,n416} ), .pin( {n441,n415} ), .gout( {n526} ), .pout( {n525} ) );
	black black_23_5 ( .gin( {n446,n416} ), .pin( {n445,n415} ), .gout( {n528} ), .pout( {n527} ) );
	black black_24_5 ( .gin( {n450,n416} ), .pin( {n449,n415} ), .gout( {n530} ), .pout( {n529} ) );
	black black_25_5 ( .gin( {n454,n416} ), .pin( {n453,n415} ), .gout( {n532} ), .pout( {n531} ) );
	black black_26_5 ( .gin( {n458,n416} ), .pin( {n457,n415} ), .gout( {n534} ), .pout( {n533} ) );
	black black_27_5 ( .gin( {n462,n416} ), .pin( {n461,n415} ), .gout( {n536} ), .pout( {n535} ) );
	black black_28_5 ( .gin( {n466,n416} ), .pin( {n465,n415} ), .gout( {n538} ), .pout( {n537} ) );
	black black_29_5 ( .gin( {n470,n416} ), .pin( {n469,n415} ), .gout( {n540} ), .pout( {n539} ) );
	black black_30_5 ( .gin( {n474,n416} ), .pin( {n473,n415} ), .gout( {n542} ), .pout( {n541} ) );
	black black_31_5 ( .gin( {n478,n416} ), .pin( {n477,n415} ), .gout( {n544} ), .pout( {n543} ) );
	post_node post_node_0_6 ( .pin( {p0} ), .gin( {n482} ), .sum( {sum[0]} ) );
	post_node post_node_1_6 ( .pin( {p1} ), .gin( {n484} ), .sum( {sum[1]} ) );
	post_node post_node_2_6 ( .pin( {p2} ), .gin( {n486} ), .sum( {sum[2]} ) );
	post_node post_node_3_6 ( .pin( {p3} ), .gin( {n488} ), .sum( {sum[3]} ) );
	post_node post_node_4_6 ( .pin( {p4} ), .gin( {n490} ), .sum( {sum[4]} ) );
	post_node post_node_5_6 ( .pin( {p5} ), .gin( {n492} ), .sum( {sum[5]} ) );
	post_node post_node_6_6 ( .pin( {p6} ), .gin( {n494} ), .sum( {sum[6]} ) );
	post_node post_node_7_6 ( .pin( {p7} ), .gin( {n496} ), .sum( {sum[7]} ) );
	post_node post_node_8_6 ( .pin( {p8} ), .gin( {n498} ), .sum( {sum[8]} ) );
	post_node post_node_9_6 ( .pin( {p9} ), .gin( {n500} ), .sum( {sum[9]} ) );
	post_node post_node_10_6 ( .pin( {p10} ), .gin( {n502} ), .sum( {sum[10]} ) );
	post_node post_node_11_6 ( .pin( {p11} ), .gin( {n504} ), .sum( {sum[11]} ) );
	post_node post_node_12_6 ( .pin( {p12} ), .gin( {n506} ), .sum( {sum[12]} ) );
	post_node post_node_13_6 ( .pin( {p13} ), .gin( {n508} ), .sum( {sum[13]} ) );
	post_node post_node_14_6 ( .pin( {p14} ), .gin( {n510} ), .sum( {sum[14]} ) );
	post_node post_node_15_6 ( .pin( {p15} ), .gin( {n512} ), .sum( {sum[15]} ) );
	post_node post_node_16_6 ( .pin( {p16} ), .gin( {n514} ), .sum( {sum[16]} ) );
	post_node post_node_17_6 ( .pin( {p17} ), .gin( {n516} ), .sum( {sum[17]} ) );
	post_node post_node_18_6 ( .pin( {p18} ), .gin( {n518} ), .sum( {sum[18]} ) );
	post_node post_node_19_6 ( .pin( {p19} ), .gin( {n520} ), .sum( {sum[19]} ) );
	post_node post_node_20_6 ( .pin( {p20} ), .gin( {n522} ), .sum( {sum[20]} ) );
	post_node post_node_21_6 ( .pin( {p21} ), .gin( {n524} ), .sum( {sum[21]} ) );
	post_node post_node_22_6 ( .pin( {p22} ), .gin( {n526} ), .sum( {sum[22]} ) );
	post_node post_node_23_6 ( .pin( {p23} ), .gin( {n528} ), .sum( {sum[23]} ) );
	post_node post_node_24_6 ( .pin( {p24} ), .gin( {n530} ), .sum( {sum[24]} ) );
	post_node post_node_25_6 ( .pin( {p25} ), .gin( {n532} ), .sum( {sum[25]} ) );
	post_node post_node_26_6 ( .pin( {p26} ), .gin( {n534} ), .sum( {sum[26]} ) );
	post_node post_node_27_6 ( .pin( {p27} ), .gin( {n536} ), .sum( {sum[27]} ) );
	post_node post_node_28_6 ( .pin( {p28} ), .gin( {n538} ), .sum( {sum[28]} ) );
	post_node post_node_29_6 ( .pin( {p29} ), .gin( {n540} ), .sum( {sum[29]} ) );
	post_node post_node_30_6 ( .pin( {p30} ), .gin( {n542} ), .sum( {sum[30]} ) );
	post_node post_node_31_6 ( .pin( {p31} ), .gin( {n544} ), .sum( {sum[31]} ) );

endmodule

module pre_node(a_in, b_in, pout, gout);

    input a_in, b_in;
    output pout, gout;

    assign pout=a_in^b_in;
    assign gout=a_in&b_in;

endmodule

module fake_pre(cin, pout, gout);

    input cin;
    output pout, gout;

    assign pout=1'b0;
    assign gout=cin;

endmodule

module post_node(pin, gin, sum);

    input pin, gin;
    output sum;

    assign sum=pin^gin;

endmodule

module invis_node(pin, gin, pout, gout);

    input pin, gin;
    output pout, gout;

    assign pout=pin;
    assign gout=gin;

endmodule

module grey(gin, pin, gout);

    input[1:0] gin;
    input pin;
    output gout;

    assign gout=gin[1]|(pin&gin[0]);

endmodule

module black(gin, pin, gout, pout);

    input [1:0] gin, pin;
    output gout, pout;

    assign pout=pin[1]&pin[0];
    assign gout=gin[1]|(pin[1]&gin[0]);

endmodule

