module adder(cout, sum, a, b, cin);

	input [31:0] a, b;
	input cin;
	output [31:0] sum;
	output cout;

	wire p9, g16, p8, g2, g9, g5, g0, g18, p6, g17, p16, p4, p0, g6, g13, g21, g29, p17, g23, p2, g_lsb, g28, g25, g26, g8, g15, p11, p14, g7, g11, p13, p28, p25, g24, p23, g12, p12, p18, p19, p27, p3, p1, p24, p29, g3, g1, p22, g20, p21, g22, p7, g19, p5, p_lsb, p15, p26, p20, g30, g4, g10, p10, g27, g14, p30;
	wire n4097, n4098, n4101, n4102, n97, n98, n99, n100, n101, n102, n105, n106, n109, n110, n111, n112, n113, n114, n117, n118, n121, n122, n123, n124, n125, n126, n129, n130, n133, n134, n135, n136, n137, n138, n141, n142, n145, n146, n147, n148, n149, n150, n153, n154, n157, n158, n159, n160, n161, n162, n165, n166, n169, n170, n171, n172, n173, n174, n177, n178, n181, n182, n183, n184, n185, n186, n189, n190, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n205, n206, n209, n210, n213, n214, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n229, n230, n233, n234, n237, n238, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n4347, n253, n254, n4348, n4351, n257, n258, n4352, n261, n262, n4355, n4356, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n4367, n4368, n277, n278, n4371, n281, n282, n4372, n285, n286, n4375, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n4395, n4396, n309, n310, n4403, n4404, n313, n314, n4411, n4412, n317, n318, n4407, n4408, n321, n322, n4419, n4420, n325, n326, n4415, n4416, n329, n330, n4427, n4428, n333, n334, n4431, n4432, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n348, n4443, n357, n358, n4451, n4452, n361, n362, n4459, n4460, n365, n366, n4463, n4464, n369, n370, n4467, n4468, n373, n374, n4471, n4472, n377, n378, n381, n382, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n421, n422, n425, n426, n429, n430, n433, n434, n437, n438, n441, n442, n445, n446, n449, n450, n453, n454, n457, n458, n461, n462, n465, n466, n469, n470, n473, n474, n477, n478, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n501, n502, n500, n503, n505, n506, n507, n508, n509, n510, n504, n511, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n537, n538, n539, n540, n541, n542, n543, n544, n512, n536, n4821, n4822, n4825, n4826, n4829, n4830, n4833, n4834, n4837, n4838, n4841, n4842, n4845, n4846, n4849, n4850, n4853, n4854, n4857, n4858, n4861, n4862, n4865, n4866, n4869, n4870, n4873, n4874, n4877, n4878, n4881, n4882, n4885, n4886, n4889, n4890, n4893, n4894, n4897, n4898, n4901, n4902, n4905, n4906, n4909, n4910, n4913, n4914, n4917, n4918, n4921, n4922, n4925, n4926, n4929, n4930, n4933, n4934, n4937, n4938, n4941, n4942, n4945, n4946, n5363, n5364, n5367, n5368, n5371, n5372, n5375, n5376, n5379, n5380, n5383, n5384, n5387, n5388, n5391, n5392, n5395, n5396, n5399, n5400, n5403, n5404, n5407, n5408, n5411, n5412, n5415, n5416, n5419, n5420, n5423, n5424, n5427, n5428, n5431, n5432, n5435, n5436, n5439, n5440, n5443, n5444, n5447, n5448, n5451, n5452, n5455, n5456, n5459, n5460, n5463, n5464, n5467, n5468, n5471, n5472, n5475, n5476, n5479, n5480, n5483, n5484, n5487, n5488, n4359, n4360, n4363, n4364, n4376, n4379, n4380, n4383, n4384, n4387, n4388, n4391, n4392, n4399, n4400, n4423, n4424, n4435, n4436, n4439, n4440, n4444, n4447, n4448, n3977, n3978, n3981, n3982, n4455, n3985, n3986, n4456, n3989, n3990, n3993, n3994, n3997, n3998, n4001, n4002, n4005, n4006, n4009, n4010, n4013, n4014, n4017, n4018, n4021, n4022, n4025, n4026, n4029, n4030, n4033, n4034, n4037, n4038, n4041, n4042, n4045, n4046, n4049, n4050, n4053, n4054, n4057, n4058, n4061, n4062, n4065, n4066, n4069, n4070, n4073, n4074, n4077, n4078, n4081, n4082, n4085, n4086, n4089, n4090, n4093, n4094;

	ppa_first_pre ppa_first_pre_0_0 ( .cin( {cin} ), .pout( {p_lsb} ), .gout( {g_lsb} ) );
	ppa_pre ppa_pre_1_0 ( .a_in( {a[0]} ), .b_in( {b[0]} ), .pout( {p0} ), .gout( {g0} ) );
	ppa_pre ppa_pre_2_0 ( .a_in( {a[1]} ), .b_in( {b[1]} ), .pout( {p1} ), .gout( {g1} ) );
	ppa_pre ppa_pre_3_0 ( .a_in( {a[2]} ), .b_in( {b[2]} ), .pout( {p2} ), .gout( {g2} ) );
	ppa_pre ppa_pre_4_0 ( .a_in( {a[3]} ), .b_in( {b[3]} ), .pout( {p3} ), .gout( {g3} ) );
	ppa_pre ppa_pre_5_0 ( .a_in( {a[4]} ), .b_in( {b[4]} ), .pout( {p4} ), .gout( {g4} ) );
	ppa_pre ppa_pre_6_0 ( .a_in( {a[5]} ), .b_in( {b[5]} ), .pout( {p5} ), .gout( {g5} ) );
	ppa_pre ppa_pre_7_0 ( .a_in( {a[6]} ), .b_in( {b[6]} ), .pout( {p6} ), .gout( {g6} ) );
	ppa_pre ppa_pre_8_0 ( .a_in( {a[7]} ), .b_in( {b[7]} ), .pout( {p7} ), .gout( {g7} ) );
	ppa_pre ppa_pre_9_0 ( .a_in( {a[8]} ), .b_in( {b[8]} ), .pout( {p8} ), .gout( {g8} ) );
	ppa_pre ppa_pre_10_0 ( .a_in( {a[9]} ), .b_in( {b[9]} ), .pout( {p9} ), .gout( {g9} ) );
	ppa_pre ppa_pre_11_0 ( .a_in( {a[10]} ), .b_in( {b[10]} ), .pout( {p10} ), .gout( {g10} ) );
	ppa_pre ppa_pre_12_0 ( .a_in( {a[11]} ), .b_in( {b[11]} ), .pout( {p11} ), .gout( {g11} ) );
	ppa_pre ppa_pre_13_0 ( .a_in( {a[12]} ), .b_in( {b[12]} ), .pout( {p12} ), .gout( {g12} ) );
	ppa_pre ppa_pre_14_0 ( .a_in( {a[13]} ), .b_in( {b[13]} ), .pout( {p13} ), .gout( {g13} ) );
	ppa_pre ppa_pre_15_0 ( .a_in( {a[14]} ), .b_in( {b[14]} ), .pout( {p14} ), .gout( {g14} ) );
	ppa_pre ppa_pre_16_0 ( .a_in( {a[15]} ), .b_in( {b[15]} ), .pout( {p15} ), .gout( {g15} ) );
	ppa_pre ppa_pre_17_0 ( .a_in( {a[16]} ), .b_in( {b[16]} ), .pout( {p16} ), .gout( {g16} ) );
	ppa_pre ppa_pre_18_0 ( .a_in( {a[17]} ), .b_in( {b[17]} ), .pout( {p17} ), .gout( {g17} ) );
	ppa_pre ppa_pre_19_0 ( .a_in( {a[18]} ), .b_in( {b[18]} ), .pout( {p18} ), .gout( {g18} ) );
	ppa_pre ppa_pre_20_0 ( .a_in( {a[19]} ), .b_in( {b[19]} ), .pout( {p19} ), .gout( {g19} ) );
	ppa_pre ppa_pre_21_0 ( .a_in( {a[20]} ), .b_in( {b[20]} ), .pout( {p20} ), .gout( {g20} ) );
	ppa_pre ppa_pre_22_0 ( .a_in( {a[21]} ), .b_in( {b[21]} ), .pout( {p21} ), .gout( {g21} ) );
	ppa_pre ppa_pre_23_0 ( .a_in( {a[22]} ), .b_in( {b[22]} ), .pout( {p22} ), .gout( {g22} ) );
	ppa_pre ppa_pre_24_0 ( .a_in( {a[23]} ), .b_in( {b[23]} ), .pout( {p23} ), .gout( {g23} ) );
	ppa_pre ppa_pre_25_0 ( .a_in( {a[24]} ), .b_in( {b[24]} ), .pout( {p24} ), .gout( {g24} ) );
	ppa_pre ppa_pre_26_0 ( .a_in( {a[25]} ), .b_in( {b[25]} ), .pout( {p25} ), .gout( {g25} ) );
	ppa_pre ppa_pre_27_0 ( .a_in( {a[26]} ), .b_in( {b[26]} ), .pout( {p26} ), .gout( {g26} ) );
	ppa_pre ppa_pre_28_0 ( .a_in( {a[27]} ), .b_in( {b[27]} ), .pout( {p27} ), .gout( {g27} ) );
	ppa_pre ppa_pre_29_0 ( .a_in( {a[28]} ), .b_in( {b[28]} ), .pout( {p28} ), .gout( {g28} ) );
	ppa_pre ppa_pre_30_0 ( .a_in( {a[29]} ), .b_in( {b[29]} ), .pout( {p29} ), .gout( {g29} ) );
	ppa_pre ppa_pre_31_0 ( .a_in( {a[30]} ), .b_in( {b[30]} ), .pout( {p30} ), .gout( {g30} ) );

	ppa_post ppa_post_0_10 ( .pin( {p0} ), .gin( {n5364} ), .sum( {sum[0]} ) );
	ppa_post ppa_post_1_10 ( .pin( {p1} ), .gin( {n5368} ), .sum( {sum[1]} ) );
	ppa_post ppa_post_2_10 ( .pin( {p2} ), .gin( {n5372} ), .sum( {sum[2]} ) );
	ppa_post ppa_post_3_10 ( .pin( {p3} ), .gin( {n5376} ), .sum( {sum[3]} ) );
	ppa_post ppa_post_4_10 ( .pin( {p4} ), .gin( {n5380} ), .sum( {sum[4]} ) );
	ppa_post ppa_post_5_10 ( .pin( {p5} ), .gin( {n5384} ), .sum( {sum[5]} ) );
	ppa_post ppa_post_6_10 ( .pin( {p6} ), .gin( {n5388} ), .sum( {sum[6]} ) );
	ppa_post ppa_post_7_10 ( .pin( {p7} ), .gin( {n5392} ), .sum( {sum[7]} ) );
	ppa_post ppa_post_8_10 ( .pin( {p8} ), .gin( {n5396} ), .sum( {sum[8]} ) );
	ppa_post ppa_post_9_10 ( .pin( {p9} ), .gin( {n5400} ), .sum( {sum[9]} ) );
	ppa_post ppa_post_10_10 ( .pin( {p10} ), .gin( {n5404} ), .sum( {sum[10]} ) );
	ppa_post ppa_post_11_10 ( .pin( {p11} ), .gin( {n5408} ), .sum( {sum[11]} ) );
	ppa_post ppa_post_12_10 ( .pin( {p12} ), .gin( {n5412} ), .sum( {sum[12]} ) );
	ppa_post ppa_post_13_10 ( .pin( {p13} ), .gin( {n5416} ), .sum( {sum[13]} ) );
	ppa_post ppa_post_14_10 ( .pin( {p14} ), .gin( {n5420} ), .sum( {sum[14]} ) );
	ppa_post ppa_post_15_10 ( .pin( {p15} ), .gin( {n5424} ), .sum( {sum[15]} ) );
	ppa_post ppa_post_16_10 ( .pin( {p16} ), .gin( {n5428} ), .sum( {sum[16]} ) );
	ppa_post ppa_post_17_10 ( .pin( {p17} ), .gin( {n5432} ), .sum( {sum[17]} ) );
	ppa_post ppa_post_18_10 ( .pin( {p18} ), .gin( {n5436} ), .sum( {sum[18]} ) );
	ppa_post ppa_post_19_10 ( .pin( {p19} ), .gin( {n5440} ), .sum( {sum[19]} ) );
	ppa_post ppa_post_20_10 ( .pin( {p20} ), .gin( {n5444} ), .sum( {sum[20]} ) );
	ppa_post ppa_post_21_10 ( .pin( {p21} ), .gin( {n5448} ), .sum( {sum[21]} ) );
	ppa_post ppa_post_22_10 ( .pin( {p22} ), .gin( {n5452} ), .sum( {sum[22]} ) );
	ppa_post ppa_post_23_10 ( .pin( {p23} ), .gin( {n5456} ), .sum( {sum[23]} ) );
	ppa_post ppa_post_24_10 ( .pin( {p24} ), .gin( {n5460} ), .sum( {sum[24]} ) );
	ppa_post ppa_post_25_10 ( .pin( {p25} ), .gin( {n5464} ), .sum( {sum[25]} ) );
	ppa_post ppa_post_26_10 ( .pin( {p26} ), .gin( {n5468} ), .sum( {sum[26]} ) );
	ppa_post ppa_post_27_10 ( .pin( {p27} ), .gin( {n5472} ), .sum( {sum[27]} ) );
	ppa_post ppa_post_28_10 ( .pin( {p28} ), .gin( {n5476} ), .sum( {sum[28]} ) );
	ppa_post ppa_post_29_10 ( .pin( {p29} ), .gin( {n5480} ), .sum( {sum[29]} ) );
	ppa_post ppa_post_30_10 ( .pin( {p30} ), .gin( {n5484} ), .sum( {sum[30]} ) );
	ppa_post ppa_post_31_10 ( .pin( {p31} ), .gin( {n5488} ), .sum( {sum[31]} ) );

	ppa_pre ppa_pre_cout ( .a_in( a[31] ), .b_in( b[31] ), .pout ( p31 ), .gout ( g31 ) );
	ppa_grey ppa_grey_cout ( .gin ( {g31,n5488} ), .pin ( p31 ), .gout ( cout ) );


    assign n97=p_lsb;
    assign n98=g_lsb;
	ppa_black ppa_black_1_1 ( .gin( {g0,g_lsb} ), .pin( {p0,p_lsb} ), .gout( {n100} ), .pout( {n99} ) );
    assign n101=p1;
    assign n102=g1;
	ppa_black ppa_black_3_1 ( .gin( {g2,g1} ), .pin( {p2,p1} ), .gout( {n106} ), .pout( {n105} ) );
    assign n109=p3;
    assign n110=g3;
	ppa_black ppa_black_5_1 ( .gin( {g4,g3} ), .pin( {p4,p3} ), .gout( {n112} ), .pout( {n111} ) );
    assign n113=p5;
    assign n114=g5;
	ppa_black ppa_black_7_1 ( .gin( {g6,g5} ), .pin( {p6,p5} ), .gout( {n118} ), .pout( {n117} ) );
    assign n121=p7;
    assign n122=g7;
	ppa_black ppa_black_9_1 ( .gin( {g8,g7} ), .pin( {p8,p7} ), .gout( {n124} ), .pout( {n123} ) );
    assign n125=p9;
    assign n126=g9;
	ppa_black ppa_black_11_1 ( .gin( {g10,g9} ), .pin( {p10,p9} ), .gout( {n130} ), .pout( {n129} ) );
    assign n133=p11;
    assign n134=g11;
	ppa_black ppa_black_13_1 ( .gin( {g12,g11} ), .pin( {p12,p11} ), .gout( {n136} ), .pout( {n135} ) );
    assign n137=p13;
    assign n138=g13;
	ppa_black ppa_black_15_1 ( .gin( {g14,g13} ), .pin( {p14,p13} ), .gout( {n142} ), .pout( {n141} ) );
    assign n145=p15;
    assign n146=g15;
	ppa_black ppa_black_17_1 ( .gin( {g16,g15} ), .pin( {p16,p15} ), .gout( {n148} ), .pout( {n147} ) );
    assign n149=p17;
    assign n150=g17;
	ppa_black ppa_black_19_1 ( .gin( {g18,g17} ), .pin( {p18,p17} ), .gout( {n154} ), .pout( {n153} ) );
    assign n157=p19;
    assign n158=g19;
	ppa_black ppa_black_21_1 ( .gin( {g20,g19} ), .pin( {p20,p19} ), .gout( {n160} ), .pout( {n159} ) );
    assign n161=p21;
    assign n162=g21;
	ppa_black ppa_black_23_1 ( .gin( {g22,g21} ), .pin( {p22,p21} ), .gout( {n166} ), .pout( {n165} ) );
    assign n169=p23;
    assign n170=g23;
	ppa_black ppa_black_25_1 ( .gin( {g24,g23} ), .pin( {p24,p23} ), .gout( {n172} ), .pout( {n171} ) );
    assign n173=p25;
    assign n174=g25;
	ppa_black ppa_black_27_1 ( .gin( {g26,g25} ), .pin( {p26,p25} ), .gout( {n178} ), .pout( {n177} ) );
    assign n181=p27;
    assign n182=g27;
	ppa_black ppa_black_29_1 ( .gin( {g28,g27} ), .pin( {p28,p27} ), .gout( {n184} ), .pout( {n183} ) );
    assign n185=p29;
    assign n186=g29;
	ppa_black ppa_black_31_1 ( .gin( {g30,g29} ), .pin( {p30,p29} ), .gout( {n190} ), .pout( {n189} ) );

    assign n193=n97;
    assign n194=n98;
    assign n195=n99;
    assign n196=n100;
    assign n197=n101;
    assign n198=n102;
	ppa_black ppa_black_3_2 ( .gin( {n106,n100} ), .pin( {n105,n99} ), .gout( {n200} ), .pout( {n199} ) );
    assign n201=n109;
    assign n202=n110;
    assign n205=n111;
    assign n206=n112;
    assign n209=n113;
    assign n210=n114;
	ppa_black ppa_black_7_2 ( .gin( {n118,n112} ), .pin( {n117,n111} ), .gout( {n214} ), .pout( {n213} ) );
    assign n217=n121;
    assign n218=n122;
    assign n219=n123;
    assign n220=n124;
    assign n221=n125;
    assign n222=n126;
	ppa_black ppa_black_11_2 ( .gin( {n130,n124} ), .pin( {n129,n123} ), .gout( {n224} ), .pout( {n223} ) );
    assign n225=n133;
    assign n226=n134;
    assign n229=n135;
    assign n230=n136;
    assign n233=n137;
    assign n234=n138;
	ppa_black ppa_black_15_2 ( .gin( {n142,n136} ), .pin( {n141,n135} ), .gout( {n238} ), .pout( {n237} ) );
    assign n241=n145;
    assign n242=n146;
    assign n243=n147;
    assign n244=n148;
    assign n245=n149;
    assign n246=n150;
	ppa_black ppa_black_19_2 ( .gin( {n154,n148} ), .pin( {n153,n147} ), .gout( {n248} ), .pout( {n247} ) );
    assign n249=n157;
    assign n250=n158;
    assign n253=n159;
    assign n254=n160;
    assign n257=n161;
    assign n258=n162;
	ppa_black ppa_black_23_2 ( .gin( {n166,n160} ), .pin( {n165,n159} ), .gout( {n262} ), .pout( {n261} ) );
    assign n265=n169;
    assign n266=n170;
    assign n267=n171;
    assign n268=n172;
    assign n269=n173;
    assign n270=n174;
	ppa_black ppa_black_27_2 ( .gin( {n178,n172} ), .pin( {n177,n171} ), .gout( {n272} ), .pout( {n271} ) );
    assign n273=n181;
    assign n274=n182;
    assign n277=n183;
    assign n278=n184;
    assign n281=n185;
    assign n282=n186;
	ppa_black ppa_black_31_2 ( .gin( {n190,n184} ), .pin( {n189,n183} ), .gout( {n286} ), .pout( {n285} ) );

    assign n289=n193;
    assign n290=n194;
    assign n291=n195;
    assign n292=n196;
    assign n293=n197;
    assign n294=n198;
    assign n295=n199;
    assign n296=n200;
    assign n297=n201;
    assign n298=n202;
    assign n299=n205;
    assign n300=n206;
    assign n301=n209;
    assign n302=n210;
	ppa_black ppa_black_7_3 ( .gin( {n214,n200} ), .pin( {n213,n199} ), .gout( {n304} ), .pout( {n303} ) );
    assign n305=n217;
    assign n306=n218;
    assign n309=n219;
    assign n310=n220;
    assign n313=n221;
    assign n314=n222;
    assign n317=n223;
    assign n318=n224;
    assign n321=n225;
    assign n322=n226;
    assign n325=n229;
    assign n326=n230;
    assign n329=n233;
    assign n330=n234;
	ppa_black ppa_black_15_3 ( .gin( {n238,n224} ), .pin( {n237,n223} ), .gout( {n334} ), .pout( {n333} ) );
    assign n337=n241;
    assign n338=n242;
    assign n339=n243;
    assign n340=n244;
    assign n341=n245;
    assign n342=n246;
    assign n343=n247;
    assign n344=n248;
    assign n345=n249;
    assign n346=n250;
    assign n347=n253;
    assign n348=n254;
    assign n349=n257;
    assign n350=n258;
	ppa_black ppa_black_23_3 ( .gin( {n262,n248} ), .pin( {n261,n247} ), .gout( {n352} ), .pout( {n351} ) );
    assign n353=n265;
    assign n354=n266;
    assign n357=n267;
    assign n358=n268;
    assign n361=n269;
    assign n362=n270;
    assign n365=n271;
    assign n366=n272;
    assign n369=n273;
    assign n370=n274;
    assign n373=n277;
    assign n374=n278;
    assign n377=n281;
    assign n378=n282;
	ppa_black ppa_black_31_3 ( .gin( {n286,n272} ), .pin( {n285,n271} ), .gout( {n382} ), .pout( {n381} ) );

    assign n385=n289;
    assign n386=n290;
    assign n387=n291;
    assign n388=n292;
    assign n389=n293;
    assign n390=n294;
    assign n391=n295;
    assign n392=n296;
    assign n393=n297;
    assign n394=n298;
    assign n395=n299;
    assign n396=n300;
    assign n397=n301;
    assign n398=n302;
    assign n399=n303;
    assign n400=n304;
    assign n401=n305;
    assign n402=n306;
    assign n403=n309;
    assign n404=n310;
    assign n405=n313;
    assign n406=n314;
    assign n407=n317;
    assign n408=n318;
    assign n409=n321;
    assign n410=n322;
    assign n411=n325;
    assign n412=n326;
    assign n413=n329;
    assign n414=n330;
	ppa_black ppa_black_15_4 ( .gin( {n334,n304} ), .pin( {n333,n303} ), .gout( {n416} ), .pout( {n415} ) );
    assign n417=n337;
    assign n418=n338;
    assign n421=n339;
    assign n422=n340;
    assign n425=n341;
    assign n426=n342;
    assign n429=n343;
    assign n430=n344;
    assign n433=n345;
    assign n434=n346;
    assign n437=n347;
    assign n438=n348;
    assign n441=n349;
    assign n442=n350;
    assign n445=n351;
    assign n446=n352;
    assign n449=n353;
    assign n450=n354;
    assign n453=n357;
    assign n454=n358;
    assign n457=n361;
    assign n458=n362;
    assign n461=n365;
    assign n462=n366;
    assign n465=n369;
    assign n466=n370;
    assign n469=n373;
    assign n470=n374;
    assign n473=n377;
    assign n474=n378;
	ppa_black ppa_black_31_4 ( .gin( {n382,n352} ), .pin( {n381,n351} ), .gout( {n478} ), .pout( {n477} ) );

    assign n481=n385;
    assign n482=n386;
	buffer_node buffer_node_1_5 ( .gin( {n388} ), .pin( {n387} ), .gout( {n484} ), .pout( {n483} ) );
    assign n485=n389;
    assign n486=n390;
	buffer_node buffer_node_3_5 ( .gin( {n392} ), .pin( {n391} ), .gout( {n488} ), .pout( {n487} ) );
    assign n489=n393;
    assign n490=n394;
    assign n491=n395;
    assign n492=n396;
    assign n493=n397;
    assign n494=n398;
	buffer_node buffer_node_7_5 ( .gin( {n400} ), .pin( {n399} ), .gout( {n496} ), .pout( {n495} ) );
    assign n497=n401;
    assign n498=n402;
    assign n499=n403;
    assign n500=n404;
    assign n501=n405;
    assign n502=n406;
    assign n503=n407;
    assign n504=n408;
    assign n505=n409;
    assign n506=n410;
    assign n507=n411;
    assign n508=n412;
    assign n509=n413;
    assign n510=n414;
	buffer_node buffer_node_15_5 ( .gin( {n416} ), .pin( {n415} ), .gout( {n512} ), .pout( {n511} ) );
    assign n513=n417;
    assign n514=n418;
    assign n515=n421;
    assign n516=n422;
    assign n517=n425;
    assign n518=n426;
    assign n519=n429;
    assign n520=n430;
    assign n521=n433;
    assign n522=n434;
    assign n523=n437;
    assign n524=n438;
    assign n525=n441;
    assign n526=n442;
    assign n527=n445;
    assign n528=n446;
    assign n529=n449;
    assign n530=n450;
    assign n531=n453;
    assign n532=n454;
    assign n533=n457;
    assign n534=n458;
    assign n535=n461;
    assign n536=n462;
    assign n537=n465;
    assign n538=n466;
    assign n539=n469;
    assign n540=n470;
    assign n541=n473;
    assign n542=n474;
	ppa_black ppa_black_31_5 ( .gin( {n478,n416} ), .pin( {n477,n415} ), .gout( {n544} ), .pout( {n543} ) );

    assign n3977=n481;
    assign n3978=n482;
    assign n3981=n483;
    assign n3982=n484;
	ppa_black ppa_black_2_6 ( .gin( {n486,n484} ), .pin( {n485,n483} ), .gout( {n3986} ), .pout( {n3985} ) );
	buffer_node buffer_node_3_6 ( .gin( {n488} ), .pin( {n487} ), .gout( {n3990} ), .pout( {n3989} ) );
    assign n3993=n489;
    assign n3994=n490;
	ppa_black ppa_black_5_6 ( .gin( {n492,n488} ), .pin( {n491,n487} ), .gout( {n3998} ), .pout( {n3997} ) );
    assign n4001=n493;
    assign n4002=n494;
	buffer_node buffer_node_7_6 ( .gin( {n496} ), .pin( {n495} ), .gout( {n4006} ), .pout( {n4005} ) );
    assign n4009=n497;
    assign n4010=n498;
    assign n4013=n499;
    assign n4014=n500;
    assign n4017=n501;
    assign n4018=n502;
	ppa_black ppa_black_11_6 ( .gin( {n504,n496} ), .pin( {n503,n495} ), .gout( {n4022} ), .pout( {n4021} ) );
    assign n4025=n505;
    assign n4026=n506;
    assign n4029=n507;
    assign n4030=n508;
    assign n4033=n509;
    assign n4034=n510;
	buffer_node buffer_node_15_6 ( .gin( {n512} ), .pin( {n511} ), .gout( {n4038} ), .pout( {n4037} ) );
    assign n4041=n513;
    assign n4042=n514;
    assign n4045=n515;
    assign n4046=n516;
    assign n4049=n517;
    assign n4050=n518;
    assign n4053=n519;
    assign n4054=n520;
    assign n4057=n521;
    assign n4058=n522;
    assign n4061=n523;
    assign n4062=n524;
    assign n4065=n525;
    assign n4066=n526;
	ppa_black ppa_black_23_6 ( .gin( {n528,n512} ), .pin( {n527,n511} ), .gout( {n4070} ), .pout( {n4069} ) );
    assign n4073=n529;
    assign n4074=n530;
    assign n4077=n531;
    assign n4078=n532;
    assign n4081=n533;
    assign n4082=n534;
    assign n4085=n535;
    assign n4086=n536;
    assign n4089=n537;
    assign n4090=n538;
    assign n4093=n539;
    assign n4094=n540;
    assign n4097=n541;
    assign n4098=n542;
    assign n4101=n543;
    assign n4102=n544;

    assign n4347=n3977;
    assign n4348=n3978;
    assign n4351=n3981;
    assign n4352=n3982;
    assign n4355=n3985;
    assign n4356=n3986;
    assign n4359=n3989;
    assign n4360=n3990;
	ppa_black ppa_black_4_7 ( .gin( {n3994,n3990} ), .pin( {n3993,n3989} ), .gout( {n4364} ), .pout( {n4363} ) );
    assign n4367=n3997;
    assign n4368=n3998;
	ppa_black ppa_black_6_7 ( .gin( {n4002,n3998} ), .pin( {n4001,n3997} ), .gout( {n4372} ), .pout( {n4371} ) );
	buffer_node buffer_node_7_7 ( .gin( {n4006} ), .pin( {n4005} ), .gout( {n4376} ), .pout( {n4375} ) );
    assign n4379=n4009;
    assign n4380=n4010;
	ppa_black ppa_black_9_7 ( .gin( {n4014,n4006} ), .pin( {n4013,n4005} ), .gout( {n4384} ), .pout( {n4383} ) );
    assign n4387=n4017;
    assign n4388=n4018;
	buffer_node buffer_node_11_7 ( .gin( {n4022} ), .pin( {n4021} ), .gout( {n4392} ), .pout( {n4391} ) );
    assign n4395=n4025;
    assign n4396=n4026;
	ppa_black ppa_black_13_7 ( .gin( {n4030,n4022} ), .pin( {n4029,n4021} ), .gout( {n4400} ), .pout( {n4399} ) );
    assign n4403=n4033;
    assign n4404=n4034;
	buffer_node buffer_node_15_7 ( .gin( {n4038} ), .pin( {n4037} ), .gout( {n4408} ), .pout( {n4407} ) );
    assign n4411=n4041;
    assign n4412=n4042;
    assign n4415=n4045;
    assign n4416=n4046;
    assign n4419=n4049;
    assign n4420=n4050;
	ppa_black ppa_black_19_7 ( .gin( {n4054,n4038} ), .pin( {n4053,n4037} ), .gout( {n4424} ), .pout( {n4423} ) );
    assign n4427=n4057;
    assign n4428=n4058;
    assign n4431=n4061;
    assign n4432=n4062;
    assign n4435=n4065;
    assign n4436=n4066;
	buffer_node buffer_node_23_7 ( .gin( {n4070} ), .pin( {n4069} ), .gout( {n4440} ), .pout( {n4439} ) );
    assign n4443=n4073;
    assign n4444=n4074;
    assign n4447=n4077;
    assign n4448=n4078;
    assign n4451=n4081;
    assign n4452=n4082;
	ppa_black ppa_black_27_7 ( .gin( {n4086,n4070} ), .pin( {n4085,n4069} ), .gout( {n4456} ), .pout( {n4455} ) );
    assign n4459=n4089;
    assign n4460=n4090;
    assign n4463=n4093;
    assign n4464=n4094;
    assign n4467=n4097;
    assign n4468=n4098;
    assign n4471=n4101;
    assign n4472=n4102;

    assign n4821=n4347;
    assign n4822=n4348;
    assign n4825=n4351;
    assign n4826=n4352;
    assign n4829=n4355;
    assign n4830=n4356;
    assign n4833=n4359;
    assign n4834=n4360;
    assign n4837=n4363;
    assign n4838=n4364;
    assign n4841=n4367;
    assign n4842=n4368;
    assign n4845=n4371;
    assign n4846=n4372;
    assign n4849=n4375;
    assign n4850=n4376;
	ppa_black ppa_black_8_8 ( .gin( {n4380,n4376} ), .pin( {n4379,n4375} ), .gout( {n4854} ), .pout( {n4853} ) );
    assign n4857=n4383;
    assign n4858=n4384;
	ppa_black ppa_black_10_8 ( .gin( {n4388,n4384} ), .pin( {n4387,n4383} ), .gout( {n4862} ), .pout( {n4861} ) );
    assign n4865=n4391;
    assign n4866=n4392;
	ppa_black ppa_black_12_8 ( .gin( {n4396,n4392} ), .pin( {n4395,n4391} ), .gout( {n4870} ), .pout( {n4869} ) );
    assign n4873=n4399;
    assign n4874=n4400;
	ppa_black ppa_black_14_8 ( .gin( {n4404,n4400} ), .pin( {n4403,n4399} ), .gout( {n4878} ), .pout( {n4877} ) );
	buffer_node buffer_node_15_8 ( .gin( {n4408} ), .pin( {n4407} ), .gout( {n4882} ), .pout( {n4881} ) );
    assign n4885=n4411;
    assign n4886=n4412;
	ppa_black ppa_black_17_8 ( .gin( {n4416,n4408} ), .pin( {n4415,n4407} ), .gout( {n4890} ), .pout( {n4889} ) );
    assign n4893=n4419;
    assign n4894=n4420;
	buffer_node buffer_node_19_8 ( .gin( {n4424} ), .pin( {n4423} ), .gout( {n4898} ), .pout( {n4897} ) );
    assign n4901=n4427;
    assign n4902=n4428;
	ppa_black ppa_black_21_8 ( .gin( {n4432,n4424} ), .pin( {n4431,n4423} ), .gout( {n4906} ), .pout( {n4905} ) );
    assign n4909=n4435;
    assign n4910=n4436;
	buffer_node buffer_node_23_8 ( .gin( {n4440} ), .pin( {n4439} ), .gout( {n4914} ), .pout( {n4913} ) );
    assign n4917=n4443;
    assign n4918=n4444;
	ppa_black ppa_black_25_8 ( .gin( {n4448,n4440} ), .pin( {n4447,n4439} ), .gout( {n4922} ), .pout( {n4921} ) );
    assign n4925=n4451;
    assign n4926=n4452;
	buffer_node buffer_node_27_8 ( .gin( {n4456} ), .pin( {n4455} ), .gout( {n4930} ), .pout( {n4929} ) );
    assign n4933=n4459;
    assign n4934=n4460;
	ppa_black ppa_black_29_8 ( .gin( {n4464,n4456} ), .pin( {n4463,n4455} ), .gout( {n4938} ), .pout( {n4937} ) );
    assign n4941=n4467;
    assign n4942=n4468;
    assign n4945=n4471;
    assign n4946=n4472;

    assign n5363=n4821;
    assign n5364=n4822;
    assign n5367=n4825;
    assign n5368=n4826;
    assign n5371=n4829;
    assign n5372=n4830;
    assign n5375=n4833;
    assign n5376=n4834;
    assign n5379=n4837;
    assign n5380=n4838;
    assign n5383=n4841;
    assign n5384=n4842;
    assign n5387=n4845;
    assign n5388=n4846;
    assign n5391=n4849;
    assign n5392=n4850;
    assign n5395=n4853;
    assign n5396=n4854;
    assign n5399=n4857;
    assign n5400=n4858;
    assign n5403=n4861;
    assign n5404=n4862;
    assign n5407=n4865;
    assign n5408=n4866;
    assign n5411=n4869;
    assign n5412=n4870;
    assign n5415=n4873;
    assign n5416=n4874;
    assign n5419=n4877;
    assign n5420=n4878;
    assign n5423=n4881;
    assign n5424=n4882;
	ppa_black ppa_black_16_9 ( .gin( {n4886,n4882} ), .pin( {n4885,n4881} ), .gout( {n5428} ), .pout( {n5427} ) );
    assign n5431=n4889;
    assign n5432=n4890;
	ppa_black ppa_black_18_9 ( .gin( {n4894,n4890} ), .pin( {n4893,n4889} ), .gout( {n5436} ), .pout( {n5435} ) );
    assign n5439=n4897;
    assign n5440=n4898;
	ppa_black ppa_black_20_9 ( .gin( {n4902,n4898} ), .pin( {n4901,n4897} ), .gout( {n5444} ), .pout( {n5443} ) );
    assign n5447=n4905;
    assign n5448=n4906;
	ppa_black ppa_black_22_9 ( .gin( {n4910,n4906} ), .pin( {n4909,n4905} ), .gout( {n5452} ), .pout( {n5451} ) );
    assign n5455=n4913;
    assign n5456=n4914;
	ppa_black ppa_black_24_9 ( .gin( {n4918,n4914} ), .pin( {n4917,n4913} ), .gout( {n5460} ), .pout( {n5459} ) );
    assign n5463=n4921;
    assign n5464=n4922;
	ppa_black ppa_black_26_9 ( .gin( {n4926,n4922} ), .pin( {n4925,n4921} ), .gout( {n5468} ), .pout( {n5467} ) );
    assign n5471=n4929;
    assign n5472=n4930;
	ppa_black ppa_black_28_9 ( .gin( {n4934,n4930} ), .pin( {n4933,n4929} ), .gout( {n5476} ), .pout( {n5475} ) );
    assign n5479=n4937;
    assign n5480=n4938;
	ppa_black ppa_black_30_9 ( .gin( {n4942,n4938} ), .pin( {n4941,n4937} ), .gout( {n5484} ), .pout( {n5483} ) );
    assign n5487=n4945;
    assign n5488=n4946;


endmodule

module ppa_grey(gin, pin, gout);

    input[1:0] gin;
    input pin;
    output gout;

    assign gout=gin[1]|(pin&gin[0]);

endmodule

module buffer_node(pin, gin, pout, gout);

    input pin, gin;
    output pout, gout;

    assign pout=pin;
    assign gout=gin;

endmodule

module ppa_black(gin, pin, gout, pout);

    input [1:0] gin, pin;
    output gout, pout;

    assign pout=pin[1]&pin[0];
    assign gout=gin[1]|(pin[1]&gin[0]);

endmodule

module invis_node(pin, gin, pout, gout);

    input pin, gin;
    output pout, gout;

    assign pout=pin;
    assign gout=gin;

endmodule

module ppa_pre(a_in, b_in, pout, gout);

    input a_in, b_in;
    output pout, gout;

    assign pout=a_in^b_in;
    assign gout=a_in&b_in;

endmodule

module ppa_post(pin, gin, sum);

    input pin, gin;
    output sum;

    assign sum=pin^gin;

endmodule

module ppa_first_pre(cin, pout, gout);

    input cin;
    output pout, gout;

    assign pout=1'b0;
    assign gout=cin;

endmodule

